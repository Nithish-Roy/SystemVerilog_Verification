class transaction;
  
  rand byte a;
  
  rand byte b;
  
 	   byte c;
  
//    event my_event;
  
  function void display( string str);
    
    $display(str);
    
    //$display($time,"a = %0d b = %0d", a, b, c);
  	
  endfunction
  
endclass

