interface adder;
  
  logic [7:0] a;
  
  logic [7:0] b;
  
  logic [8:0] c;
  
endinterface
