module adder_module (input byte a, input byte b, output bit [8:0] c);
  
assign c = a + b;
  
endmodule
